mem[0] = 8'h6F;
mem[1] = 8'h00;
mem[2] = 8'h40;
mem[3] = 8'h01;
mem[4] = 8'h13;
mem[5] = 8'h00;
mem[6] = 8'h00;
mem[7] = 8'h00;
mem[8] = 8'h13;
mem[9] = 8'h00;
mem[10] = 8'h00;
mem[11] = 8'h00;
mem[12] = 8'h13;
mem[13] = 8'h00;
mem[14] = 8'h00;
mem[15] = 8'h00;
mem[16] = 8'h6F;
mem[17] = 8'h00;
mem[18] = 8'h40;
mem[19] = 8'h02;
mem[20] = 8'h93;
mem[21] = 8'h00;
mem[22] = 8'h80;
mem[23] = 8'h00;
mem[24] = 8'h93;
mem[25] = 8'hC0;
mem[26] = 8'hF0;
mem[27] = 8'hFF;
mem[28] = 8'h0B;
mem[29] = 8'hE0;
mem[30] = 8'h00;
mem[31] = 8'h06;
mem[32] = 8'h93;
mem[33] = 8'h00;
mem[34] = 8'h00;
mem[35] = 8'h00;
mem[36] = 8'h93;
mem[37] = 8'h01;
mem[38] = 8'h00;
mem[39] = 8'h00;
mem[40] = 8'h13;
mem[41] = 8'h02;
mem[42] = 8'h00;
mem[43] = 8'h00;
mem[44] = 8'h0B;
mem[45] = 8'h40;
mem[46] = 8'h00;
mem[47] = 8'h08;
mem[48] = 8'h6F;
mem[49] = 8'hF0;
mem[50] = 8'hDF;
mem[51] = 8'hFF;
mem[52] = 8'h93;
mem[53] = 8'h81;
mem[54] = 8'h11;
mem[55] = 8'h00;
mem[56] = 8'h63;
mem[57] = 8'hEA;
mem[58] = 8'h41;
mem[59] = 8'h00;
mem[60] = 8'h93;
mem[61] = 8'h01;
mem[62] = 8'h00;
mem[63] = 8'h00;
mem[64] = 8'h93;
mem[65] = 8'h80;
mem[66] = 8'h10;
mem[67] = 8'h00;
mem[68] = 8'h37;
mem[69] = 8'h11;
mem[70] = 8'h00;
mem[71] = 8'h00;
mem[72] = 8'h23;
mem[73] = 8'h20;
mem[74] = 8'h11;
mem[75] = 8'h00;
mem[76] = 8'h0B;
mem[77] = 8'h00;
mem[78] = 8'h00;
mem[79] = 8'h04;
for (i = 4016; i < 4096; i = i + 1) mem[i] = 0;